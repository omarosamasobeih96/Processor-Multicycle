LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY rom IS
	PORT( 	address : in std_logic_vector(5 downto 0);
		Ain, Bout, Cin, Cout, ALUOperation : out std_logic_vector(3 downto 0);
		rst, RamWriteEnable, SetCarry, NeedCarry, DestinationWrite, MFC, HLT, wordMode : out std_logic;
		NextRomAddressSel : out std_logic_vector(2 downto 0));
END ENTITY rom;

ARCHITECTURE arch1 OF rom IS
	--first 3 bits => src, second 3 bits => dst, rest => DataBus
	TYPE rom_data IS ARRAY(0 TO 49) OF std_logic_vector(30 DOWNTO 0);
	CONSTANT rom : rom_data := (
		 0 => "0000011111000111111110000010100",
		 1 => "0000111110110111110000000010100",
		 2 => "0000111110110111110000000110100",
		 3 => "0001011110110111110000010010100",
		 4 => "0001011110110111110000000110100",
		 5 => "0010011110110111110000000010100",
		 6 => "0010111110110111110000000010100",
		 7 => "0011011110110111110000000010100",
		 8 => "0011110001000111111110000000000",
		 9 => "0010011110110111110000000010100",
		10 => "0001011110110111110000010000100",
		11 => "0000011110110111111110010010100",
		12 => "0001111110110111111110000010100",
		13 => "0111111111111111111110000010100",
		14 => "0011111110110111111110000010100",
		15 => "0100011110110111111110000010100",
		16 => "0100111110110111111110000010100",
		17 => "0101011110110111111110000110100",
		18 => "0101111110110111111110000010100",
		19 => "0110011110110111111110000010100",
		20 => "0110111110110111111110000010100",
		21 => "0111011110110111111110000110100",
		22 => "0111111111111111111110000001100",
		23 => "0111111111111111111110000000100",
		24 => "0111111111111111111111000000100",
		25 => "1000000100010010100100011000000",
		26 => "0001101010011100001100000000000",
		27 => "1001100110011011000100101000000",
		28 => "0111111111111001010000000000100",
		29 => "1111111111111010100110001000000",
		30 => "0000000110011001001100010000100",
		31 => "0111111111111100000010000000010",
		32 => "0000000010001010100010011000000",
		33 => "0000011111111100001100000000010",
		34 => "0001101010001111111110001000000",
		35 => "0001100010001100001100000000010",
		36 => "1000000100010010100100011000000",
		37 => "0000101010001111101100001000000",
		38 => "0111111111111100001100000000010",
		39 => "0111111111111011000000000000011",
		40 => "0000000000000010100000011000011",
		41 => "0001101010000111111110001000000",
		42 => "0001100000000111111110000000011",
		43 => "1000000100010010100100011000000",
		44 => "0000101010001111101100001000011",
		45 => "1000000100010010100100011000000",
		46 => "0111111111111010001100000000001",
		47 => "1000000100010010100100011000000",
		48 => "0010010000111111101100000000000",
		49 => "0000100101000111100100000000100"
	);
BEGIN	
	wordMode <= rom(to_integer(unsigned(address)))(30);
	ALUOperation <= rom(to_integer(unsigned(address)))(29 downto 26);
	Ain <= rom(to_integer(unsigned(address)))(25 downto 22);
	Bout <= rom(to_integer(unsigned(address)))(21 downto 18);
	Cin <= rom(to_integer(unsigned(address)))(17 downto 14);
	Cout <= rom(to_integer(unsigned(address)))(13 downto 10);
	rst <= rom(to_integer(unsigned(address)))(9);
	RamWriteEnable <= rom(to_integer(unsigned(address)))(8);
	SetCarry <= rom(to_integer(unsigned(address)))(7);
	MFC <= rom(to_integer(unsigned(address)))(6);
	NeedCarry <= rom(to_integer(unsigned(address)))(5);
	DestinationWrite <= rom(to_integer(unsigned(address)))(4);
	HLT <= rom(to_integer(unsigned(address)))(3);
	NextRomAddressSel <= rom(to_integer(unsigned(address)))(2 downto 0);
END arch1;
